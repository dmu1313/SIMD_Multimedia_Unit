-------------------------------------------------------------------------------
--
-- Title       : Test
-- Design      : SIMD_Multimedia_Unit
-- Author      : Brian Eng
-- Company     : StonyBrook
--
-------------------------------------------------------------------------------
--
-- File        : c:\My_Designs\Ese_345\SIMD_Multimedia_Unit\src\Test.vhd
-- Generated   : Tue Dec  3 21:46:02 2019
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {Test} architecture {Test}}

library IEEE;
use IEEE.std_logic_1164.all;

entity Test is
	 port(
		 a : in STD_LOGIC
	     );
end Test;

--}} End of automatically maintained section

architecture Test of Test is
begin

	 -- enter your statements here --

end Test;
